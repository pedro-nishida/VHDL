ENTITY M12121ECP015 IS
PORT(
	D0, D1, D2, D3: IN BIT;			-- vARIAVEIS DE SINAL DE ENTRADA
	X: IN INTEGER RANGE 0 TO 3;	-- ENTRADA A1 E A0 EM INT
	S: OUT BIT							-- VARIAVEL DE SAIDA
);


END M12121ECP015;


ARCHITECTURE CIR OF M12121ECP015 IS
BEGIN
	WITH X SELECT
	S<=D0 WHEN 0,
		D1 WHEN 1,
		D2 WHEN 2,
		D3 WHEN 3;		
END CIR;