--PROJETO TABELA VERDADE 2
ENTITY M12121ECP015 IS
PORT(
	VET: IN INTEGER RANGE 0 TO 15; 
	S1, S2: OUT BIT
);


END M12121ECP015;


ARCHITECTURE CIR OF M12121ECP015 IS
	SIGNAL AUX:BIT_VECTOR (1 DOWNTO 0);--AUXILIAR PARA ENDEREÇAR S1 E S2
BEGIN
	WITH VET SELECT
		AUX<="10" WHEN 0,
			  "00" WHEN 1,
			  "01" WHEN 2,
			  "11" WHEN 3,
			  "01" WHEN 4,
			  "00" WHEN 5,
			  "01" WHEN 6,
			  "10" WHEN 7,
			  "10" WHEN 8,
			  "01" WHEN 9,
			  "10" WHEN 10,
			  "10" WHEN 11,
			  "10" WHEN 12,
			  "11" WHEN 13,
			  "00" WHEN 14,
			  "10" WHEN 15;
			-- ATENÇÃO ASPAS SIMPLES IMPLICA EM BIT ENQUANTO ASPAS DUPLAS IMPLICA EM VETOR
	
	-- ALOCAR QUAL INDEX DO VETOR É REFERENTE A SAIDA DESEJADA
	S1<= AUX(1);
	S2<= AUX(0);
END CIR;